


`include "/proj/repo/user/vaibhavb/ai_i2s_rtl/ai_i2s_top.sv"
`include "/proj/repo/user/vaibhavb/ai_i2s_rtl/ai_i2s_testbench.sv"                  
